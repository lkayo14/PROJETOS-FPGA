ENTITY DECODIFICADOR_7SEG IS
PORT ( DISPLAY: OUT BIT_VECTOR(6 DOWNTO 0);
DEC: IN INTEGER RANGE 0 TO 7);
END DECODIFICADOR_7SEG;

ARCHITECTURE ONE OF DECODIFICADOR_7SEG IS 
BEGIN
WITH DEC SELECT
	DISPLAY <= "0011000" WHEN 0,
		        "1001111" WHEN 1,
				  "1100000" WHEN 2,
				  "0100100" WHEN 3,
				  "0010010" WHEN 4,
				  "1110000" WHEN 5,
				  "1001100" WHEN 6,
				  "0000110" WHEN 7;
END ONE;
				  
