ENTITY COMUTADOR IS
PORT(CLK, P, B: IN BIT;
K1,K2,K3: OUT BIT;
DISPLAY_0: OUT BIT_VECTOR(6 DOWNTO 0));

END COMUTADOR;

ARCHITECTURE ONE OF COMUTADOR IS

SIGNAL AUX:BIT;

SIGNAL AUX_1: INTEGER RANGE 0 TO 7;



COMPONENT DIV_CLK IS
PORT (IN_CLK: IN BIT;
OUT_CLK: OUT BIT);
END COMPONENT;


COMPONENT FSM_1 IS
PORT (IN_CLK, S1, S2: IN BIT;
C1, C2, C3: OUT BIT;
DEC: OUT INTEGER RANGE 0 TO 7);
END COMPONENT;


COMPONENT DECODIFICADOR_7SEG IS
PORT ( DISPLAY: OUT BIT_VECTOR(6 DOWNTO 0);
IN_DEC: IN INTEGER RANGE 0 TO 7);
END COMPONENT;


BEGIN
	
	CHIP1: DIV_CLK PORT MAP(IN_CLK=>CLK, OUT_CLK=>AUX);
	
	CHIP2: FSM_1 PORT MAP(IN_CLK=>AUX,S1=>P,S2=>B,C1=>K1,C2=>K2,C3=>K3, DEC=>AUX_1);
	
	CHIP3: DECODIFICADOR_7SEG PORT MAP(DISPLAY=>DISPLAY_0,IN_DEC=>AUX_1);
	
	
END ONE;

ENTITY DIV_CLK IS
PORT ( IN_CLK: IN BIT;
OUT_CLK : OUT BIT);
END DIV_CLK;

ARCHITECTURE ONE OF DIV_CLK IS
SIGNAL X: BIT;
SIGNAL Y: INTEGER RANGE 0 TO 4 :=0;

BEGIN 
PROCESS (IN_CLK)
BEGIN
IF (IN_CLK'EVENT)AND(IN_CLK='1') THEN
  IF Y=4 THEN
  Y<=0;
  X<=NOT X;
  ELSE
  Y<= Y+1;
  END IF;
END IF;
END PROCESS;
OUT_CLK<= X;
END ONE;


ENTITY FSM_1 IS
PORT (S1,S2, IN_CLK : IN BIT;
C1, C2, C3 : OUT BIT;
DEC: OUT INTEGER RANGE 0 TO 7);
END FSM_1;

ARCHITECTURE ONE OF FSM_1 IS
TYPE STATE IS (GP, H1, GB, H5, H2, PA, H4, H3);
SIGNAL AUX : STATE;
BEGIN
PROCESS (IN_CLK)
BEGIN
IF (IN_CLK'EVENT)AND(IN_CLK='1')THEN
       CASE AUX IS 
		 WHEN GP =>
		 IF (S1='0'AND S2='1') THEN
		 AUX<=H1;
		 ELSIF (S1='0'AND S2='0') THEN
		 AUX<=H4;
		 ELSE
		 AUX<=GP;
		 END IF;
		 
		 WHEN H1 =>
		 AUX<= GB;
		 
		 WHEN GB =>
		 IF (S1='1') THEN
		 AUX<=H5;
       ELSIF (S1='0'AND S2='0') THEN
		 AUX<=H2;
		 ELSE
		 AUX<=GB;
		 END IF;
		 
		 WHEN H2 =>
		 AUX<= PA;
		 
		 WHEN H5 =>
		 AUX<= GP;
		 
		 WHEN H4 =>
		 AUX<= PA;
		 
		 WHEN PA =>
		 IF (S1='1') THEN
		 AUX<=H3;
       ELSE 
		 AUX<=PA;
		 END IF;
		 
		 WHEN H3 =>
		 AUX<= GP;
		 
		END CASE;
		END IF;
END PROCESS;
	
	
WITH AUX SELECT
	C1<= '1' WHEN GP,
		  '1' WHEN H1,
		  '1' WHEN H4,
		  '0' WHEN OTHERS;

WITH AUX SELECT
	C2<= '1' WHEN GB,
		  '1' WHEN H2,
		  '1' WHEN H5,
		  '0' WHEN OTHERS;		  
		  
WITH AUX SELECT
	C3<= '1' WHEN GP,
		  '1' WHEN H1,
		  '1' WHEN H4,
		  '0' WHEN OTHERS;	
	
WITH AUX SELECT
	DEC<= 0 WHEN GP,
		   1 WHEN H1,
		   2 WHEN GB,
		   3 WHEN H5,
			4 WHEN H2,
		   5 WHEN PA,
			6 WHEN H4,
			7 WHEN H3;
	
		 
END ONE;


ENTITY DECODIFICADOR_7SEG IS
PORT ( DISPLAY: OUT BIT_VECTOR(6 DOWNTO 0);
IN_DEC: IN INTEGER RANGE 0 TO 7);
END DECODIFICADOR_7SEG;

ARCHITECTURE ONE OF DECODIFICADOR_7SEG IS 
BEGIN
WITH IN_DEC SELECT
	DISPLAY <= "0011000" WHEN 0,
		        "1001111" WHEN 1,
				  "1100000" WHEN 2,
				  "0100100" WHEN 3,
				  "0010010" WHEN 4,
				  "1110000" WHEN 5,
				  "1001100" WHEN 6,
				  "0000110" WHEN 7;
END ONE;
				  

